module alu(
    input [15:0] AR,
    input [15:0] AC_in,
    input [7:0] INPR,
    output reg E,
    output [15:0] AC_out,
);

endmodule