module cu_PC(
    
);


endmodule