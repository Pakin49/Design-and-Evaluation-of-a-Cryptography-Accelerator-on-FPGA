module alu(
    input [3:0] Selector
    input [15:0] DR,
    input [15:0] AC_in,
    input [7:0] INPR,
    output reg E,
    output [15:0] AC,
);
assign 

endmodule