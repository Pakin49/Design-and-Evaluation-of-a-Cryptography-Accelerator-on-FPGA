module data_bus(

);

endmodule