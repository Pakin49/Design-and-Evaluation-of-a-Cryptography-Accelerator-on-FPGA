module cpu;
    `include cpu.sv
    `include alu.sv
    my_register AC(
        
    );

endmodule