module main;
    my_register AC(

    );
endmodule